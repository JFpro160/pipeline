module eqcmp #(parameter WIDTH = 8) (
    input wire [WIDTH - 1:0] a, b,
    output wire y
);
    assign y = (a == b);
endmodule